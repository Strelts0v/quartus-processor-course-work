registerMux_inst : registerMux PORT MAP (
		data0x	 => data0x_sig,
		data10x	 => data10x_sig,
		data11x	 => data11x_sig,
		data12x	 => data12x_sig,
		data13x	 => data13x_sig,
		data14x	 => data14x_sig,
		data15x	 => data15x_sig,
		data16x	 => data16x_sig,
		data17x	 => data17x_sig,
		data18x	 => data18x_sig,
		data19x	 => data19x_sig,
		data1x	 => data1x_sig,
		data20x	 => data20x_sig,
		data21x	 => data21x_sig,
		data22x	 => data22x_sig,
		data23x	 => data23x_sig,
		data24x	 => data24x_sig,
		data25x	 => data25x_sig,
		data26x	 => data26x_sig,
		data27x	 => data27x_sig,
		data2x	 => data2x_sig,
		data3x	 => data3x_sig,
		data4x	 => data4x_sig,
		data5x	 => data5x_sig,
		data6x	 => data6x_sig,
		data7x	 => data7x_sig,
		data8x	 => data8x_sig,
		data9x	 => data9x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
