address_invertor_inst : address_invertor PORT MAP (
		data	 => data_sig,
		result	 => result_sig
	);
