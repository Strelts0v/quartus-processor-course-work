lpm_add_sub0_inst : lpm_add_sub0 PORT MAP (
		dataa	 => dataa_sig,
		overflow	 => overflow_sig,
		result	 => result_sig
	);
