stack_register_inst : stack_register PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
