ab_comparator_inst : ab_comparator PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AeB	 => AeB_sig,
		AgB	 => AgB_sig,
		AlB	 => AlB_sig
	);
