lpm_add_sub3_inst : lpm_add_sub3 PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
