lpm_mux1_inst : lpm_mux1 PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
