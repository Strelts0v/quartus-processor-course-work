stack_pointer_register_inst : stack_pointer_register PORT MAP (
		aset	 => aset_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
