stack_push_counter_inst : stack_push_counter PORT MAP (
		dataa	 => dataa_sig,
		overflow	 => overflow_sig,
		result	 => result_sig
	);
