stack_address_sub_inst : stack_address_sub PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
