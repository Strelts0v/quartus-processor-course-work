lpm_add_sub2_inst : lpm_add_sub2 PORT MAP (
		dataa	 => dataa_sig,
		overflow	 => overflow_sig,
		result	 => result_sig
	);
