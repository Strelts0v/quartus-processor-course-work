ALU_ADD_inst : ALU_ADD PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		cout	 => cout_sig,
		overflow	 => overflow_sig,
		result	 => result_sig
	);
