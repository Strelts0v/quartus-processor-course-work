stack_pop_counter_inst : stack_pop_counter PORT MAP (
		dataa	 => dataa_sig,
		overflow	 => overflow_sig,
		result	 => result_sig
	);
