lpm_dff2_inst : lpm_dff2 PORT MAP (
		aset	 => aset_sig,
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
