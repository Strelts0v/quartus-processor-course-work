lpm_clshift1_inst : lpm_clshift1 PORT MAP (
		data	 => data_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
